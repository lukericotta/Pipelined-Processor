module CacheDecoder_7_128(input [6:0] RegId, input WriteReg, output [127:0] Wordline);

assign Wordline = (WriteReg == 1'b1)  ? (
		  (RegId == 7'd0) ? 128'h00000000000000000000000000000001 :
		  (RegId == 7'd1) ? 128'h00000000000000000000000000000002 :
		  (RegId == 7'd2) ? 128'h00000000000000000000000000000004 :
		  (RegId == 7'd3) ? 128'h00000000000000000000000000000008 :
		  (RegId == 7'd4) ? 128'h00000000000000000000000000000010 :
		  (RegId == 7'd5) ? 128'h00000000000000000000000000000020 :
		  (RegId == 7'd6) ? 128'h00000000000000000000000000000040 :
		  (RegId == 7'd7) ? 128'h00000000000000000000000000000080 :
		  (RegId == 7'd8) ? 128'h00000000000000000000000000000100 :
		  (RegId == 7'd9) ? 128'h00000000000000000000000000000200 :
		  (RegId == 7'd10) ? 128'h00000000000000000000000000000400 :
		  (RegId == 7'd11) ? 128'h00000000000000000000000000000800 :
		  (RegId == 7'd12) ? 128'h00000000000000000000000000001000 :
		  (RegId == 7'd13) ? 128'h00000000000000000000000000002000 :
		  (RegId == 7'd14) ? 128'h00000000000000000000000000004000 :
		  (RegId == 7'd15) ? 128'h00000000000000000000000000008000 :
		  (RegId == 7'd16) ? 128'h00000000000000000000000000010000 :
		  (RegId == 7'd17) ? 128'h00000000000000000000000000020000 :
		  (RegId == 7'd18) ? 128'h00000000000000000000000000040000 :
		  (RegId == 7'd19) ? 128'h00000000000000000000000000080000 :
		  (RegId == 7'd20) ? 128'h00000000000000000000000000100000 :
		  (RegId == 7'd21) ? 128'h00000000000000000000000000200000 :
		  (RegId == 7'd22) ? 128'h00000000000000000000000000400000 :
		  (RegId == 7'd23) ? 128'h00000000000000000000000000800000 :
		  (RegId == 7'd24) ? 128'h00000000000000000000000001000000 :
		  (RegId == 7'd25) ? 128'h00000000000000000000000002000000 :
		  (RegId == 7'd26) ? 128'h00000000000000000000000004000000 :
		  (RegId == 7'd27) ? 128'h00000000000000000000000008000000 :
		  (RegId == 7'd28) ? 128'h00000000000000000000000010000000 :
		  (RegId == 7'd29) ? 128'h00000000000000000000000020000000 :
		  (RegId == 7'd30) ? 128'h00000000000000000000000040000000 :
		  (RegId == 7'd31) ? 128'h00000000000000000000000080000000 :
		  (RegId == 7'd32) ? 128'h00000000000000000000000100000000 :
		  (RegId == 7'd33) ? 128'h00000000000000000000000200000000 :
		  (RegId == 7'd34) ? 128'h00000000000000000000000400000000 :
		  (RegId == 7'd35) ? 128'h00000000000000000000000800000000 :
		  (RegId == 7'd36) ? 128'h00000000000000000000001000000000 :
		  (RegId == 7'd37) ? 128'h00000000000000000000002000000000 :
		  (RegId == 7'd38) ? 128'h00000000000000000000004000000000 :
		  (RegId == 7'd39) ? 128'h00000000000000000000008000000000 :
		  (RegId == 7'd40) ? 128'h00000000000000000000010000000000 :
		  (RegId == 7'd41) ? 128'h00000000000000000000020000000000 :
		  (RegId == 7'd42) ? 128'h00000000000000000000040000000000 :
		  (RegId == 7'd43) ? 128'h00000000000000000000080000000000 :
		  (RegId == 7'd44) ? 128'h00000000000000000000100000000000 :
		  (RegId == 7'd45) ? 128'h00000000000000000000200000000000 :
		  (RegId == 7'd46) ? 128'h00000000000000000000400000000000 :
		  (RegId == 7'd47) ? 128'h00000000000000000000800000000000 :
		  (RegId == 7'd48) ? 128'h00000000000000000001000000000000 :
		  (RegId == 7'd49) ? 128'h00000000000000000002000000000000 :
		  (RegId == 7'd50) ? 128'h00000000000000000004000000000000 :
		  (RegId == 7'd51) ? 128'h00000000000000000008000000000000 :
		  (RegId == 7'd52) ? 128'h00000000000000000010000000000000 :
		  (RegId == 7'd53) ? 128'h00000000000000000020000000000000 :
		  (RegId == 7'd54) ? 128'h00000000000000000040000000000000 :
		  (RegId == 7'd55) ? 128'h00000000000000000080000000000000 :
		  (RegId == 7'd56) ? 128'h00000000000000000100000000000000 :
		  (RegId == 7'd57) ? 128'h00000000000000000200000000000000 :
		  (RegId == 7'd58) ? 128'h00000000000000000400000000000000 :
		  (RegId == 7'd59) ? 128'h00000000000000000800000000000000 :
		  (RegId == 7'd60) ? 128'h00000000000000001000000000000000 :
		  (RegId == 7'd61) ? 128'h00000000000000002000000000000000 :
		  (RegId == 7'd62) ? 128'h00000000000000004000000000000000 :
		  (RegId == 7'd63) ? 128'h00000000000000008000000000000000 :
		  (RegId == 7'd64) ? 128'h00000000000000010000000000000000 :
		  (RegId == 7'd65) ? 128'h00000000000000020000000000000000 :
		  (RegId == 7'd66) ? 128'h00000000000000040000000000000000 :
		  (RegId == 7'd67) ? 128'h00000000000000080000000000000000 :
		  (RegId == 7'd68) ? 128'h00000000000000100000000000000000 :
		  (RegId == 7'd69) ? 128'h00000000000000200000000000000000 :
		  (RegId == 7'd70) ? 128'h00000000000000400000000000000000 :
		  (RegId == 7'd71) ? 128'h00000000000000800000000000000000 :
		  (RegId == 7'd72) ? 128'h00000000000001000000000000000000 :
		  (RegId == 7'd73) ? 128'h00000000000002000000000000000000 :
		  (RegId == 7'd74) ? 128'h00000000000004000000000000000000 :
		  (RegId == 7'd75) ? 128'h00000000000008000000000000000000 :
		  (RegId == 7'd76) ? 128'h00000000000010000000000000000000 :
		  (RegId == 7'd77) ? 128'h00000000000020000000000000000000 :
		  (RegId == 7'd78) ? 128'h00000000000040000000000000000000 :
		  (RegId == 7'd79) ? 128'h00000000000080000000000000000000 :
		  (RegId == 7'd80) ? 128'h00000000000100000000000000000000 :
		  (RegId == 7'd81) ? 128'h00000000000200000000000000000000 :
		  (RegId == 7'd82) ? 128'h00000000000400000000000000000000 :
		  (RegId == 7'd83) ? 128'h00000000000800000000000000000000 :
		  (RegId == 7'd84) ? 128'h00000000001000000000000000000000 :
		  (RegId == 7'd85) ? 128'h00000000002000000000000000000000 :
		  (RegId == 7'd86) ? 128'h00000000004000000000000000000000 :
		  (RegId == 7'd87) ? 128'h00000000008000000000000000000000 :
		  (RegId == 7'd88) ? 128'h00000000010000000000000000000000 :
		  (RegId == 7'd89) ? 128'h00000000020000000000000000000000 :
		  (RegId == 7'd90) ? 128'h00000000040000000000000000000000 :
		  (RegId == 7'd91) ? 128'h00000000080000000000000000000000 :
		  (RegId == 7'd92) ? 128'h00000000100000000000000000000000 :
		  (RegId == 7'd93) ? 128'h00000000200000000000000000000000 :
		  (RegId == 7'd94) ? 128'h00000000400000000000000000000000 :
		  (RegId == 7'd95) ? 128'h00000000800000000000000000000000 :
		  (RegId == 7'd96) ? 128'h00000001000000000000000000000000 :
		  (RegId == 7'd97) ? 128'h00000002000000000000000000000000 :
		  (RegId == 7'd98) ? 128'h00000004000000000000000000000000 :
		  (RegId == 7'd99) ? 128'h00000008000000000000000000000000 :
		  (RegId == 7'd100) ? 128'h00000010000000000000000000000000 :
		  (RegId == 7'd101) ? 128'h00000020000000000000000000000000 :
		  (RegId == 7'd102) ? 128'h00000040000000000000000000000000 :
		  (RegId == 7'd103) ? 128'h00000080000000000000000000000000 :
		  (RegId == 7'd104) ? 128'h00000100000000000000000000000000 :
		  (RegId == 7'd105) ? 128'h00000200000000000000000000000000 :
		  (RegId == 7'd106) ? 128'h00000400000000000000000000000000 :
		  (RegId == 7'd107) ? 128'h00000800000000000000000000000000 :
		  (RegId == 7'd108) ? 128'h00001000000000000000000000000000 :
		  (RegId == 7'd109) ? 128'h00002000000000000000000000000000 :
		  (RegId == 7'd110) ? 128'h00004000000000000000000000000000 :
		  (RegId == 7'd111) ? 128'h00008000000000000000000000000000 :
		  (RegId == 7'd112) ? 128'h00010000000000000000000000000000 :
		  (RegId == 7'd113) ? 128'h00020000000000000000000000000000 :
		  (RegId == 7'd114) ? 128'h00040000000000000000000000000000 :
		  (RegId == 7'd115) ? 128'h00080000000000000000000000000000 :
		  (RegId == 7'd116) ? 128'h00100000000000000000000000000000 :
		  (RegId == 7'd117) ? 128'h00200000000000000000000000000000 :
		  (RegId == 7'd118) ? 128'h00400000000000000000000000000000 :
		  (RegId == 7'd119) ? 128'h00800000000000000000000000000000 :
		  (RegId == 7'd120) ? 128'h01000000000000000000000000000000 :
		  (RegId == 7'd121) ? 128'h02000000000000000000000000000000 :
		  (RegId == 7'd122) ? 128'h04000000000000000000000000000000 :
		  (RegId == 7'd123) ? 128'h08000000000000000000000000000000 :
		  (RegId == 7'd124) ? 128'h10000000000000000000000000000000 :
		  (RegId == 7'd125) ? 128'h20000000000000000000000000000000 :
		  (RegId == 7'd126) ? 128'h40000000000000000000000000000000 :
		  (RegId == 7'd127) ? 128'h80000000000000000000000000000000 :
					128'h00000000000000000000000000000000) 
						: 128'h00000000000000000000000000000000;

endmodule
